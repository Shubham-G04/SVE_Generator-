module generate2 (
    input wire clk,
    input wire rst,
    input wire [8-1:0] a,
    input wire [8-1:0] b,
    output wire [8-1:0] y
);

// DUT logic here

endmodule
